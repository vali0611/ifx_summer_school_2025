/******************************************************************************
 * (C) Copyright 2020 All Rights Reserved
 *
 * MODULE:
 * DEVICE:
 * PROJECT:
 * AUTHOR:
 * DATE:
 * FILE:
 * REVISION:
 *
 * FILE DESCRIPTION:
 *
 *******************************************************************************/

`timescale 1ns/100ps

package ifx_dig_data_bus_uvc_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ifx_dig_data_bus_uvc_typedef.svh"
  `include "ifx_dig_data_bus_uvc_config.svh"
  // TODO: Include data bus uvc files

endpackage
