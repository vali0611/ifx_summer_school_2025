package ifx_dig_regblock_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
   `include "ifx_dig_defines.svh"

  // TODO: Include regblock files
  `include "ifx_dig_field.svh"
  `include "ifx_dig_registers.svh"
  `include "ifx_dig_regblock.svh"

endpackage
