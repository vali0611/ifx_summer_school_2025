/******************************************************************************
 * (C) Copyright 2019 All Rights Reserved
 *
 * MODULE:
 * DEVICE:
 * PROJECT:
 * AUTHOR:
 * DATE:
 * FILE:
 * REVISION:
 *
 * FILE DESCRIPTION:
 *
 *******************************************************************************/

package ifx_dig_pkg;

  //=========================================================================
  // UVM and DEFINES.
  //-------------------------------------------------------------------------
  //=========================================================================
  import uvm_pkg::*;
  `include  "uvm_macros.svh"

  `include "ifx_dig_defines.svh"

  //=========================================================================
  // TODO: import the UVC packages
  //-------------------------------------------------------------------------
  import ifx_dig_regblock_pkg::*;

  //=========================================================================
  // TODO: Include Environment files (env, scoreboard, sequencer, types, config)
  //-------------------------------------------------------------------------
  //=========================================================================


endpackage
