/******************************************************************************
 * (C) Copyright 2020 All Rights Reserved
 *
 * MODULE:
 * DEVICE:
 * PROJECT:
 * AUTHOR:
 * DATE:
 * FILE:
 * REVISION:
 *
 * FILE DESCRIPTION:
 *
 *******************************************************************************/
 
typedef enum int {READ=0, WRITE=1, INVALID_READ=3, INVALID_WRITE=4} access_type_t;
typedef enum int {ADDR_INVALID=1, ADDR_VALID=0} address_validity_t;